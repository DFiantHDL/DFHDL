`default_nettype none
`timescale 1ns/1ps
`include "Cipher_defs.vh"

module mixColumns(
  state,
  o
);
  `include "dfhdl_defs.vh"
  `include "Cipher_defs.vh"
  input  wire  [7:0] state [0:3] [0:3];
  output wire [7:0] o [0:3] [0:3];
  wire [7:0] o_part_mulByte_0_inst_rhs;
  wire [7:0] o_part_mulByte_0_inst_o;
  wire [7:0] o_part_mulByte_1_inst_rhs;
  wire [7:0] o_part_mulByte_1_inst_o;
  wire [7:0] o_part_mulByte_2_inst_rhs;
  wire [7:0] o_part_mulByte_2_inst_o;
  wire [7:0] mulByte_2_inst_00_rhs;
  wire [7:0] mulByte_2_inst_00_o;
  wire [7:0] mulByte_2_inst_01_rhs;
  wire [7:0] mulByte_2_inst_01_o;
  wire [7:0] mulByte_0_inst_00_rhs;
  wire [7:0] mulByte_0_inst_00_o;
  wire [7:0] mulByte_1_inst_00_rhs;
  wire [7:0] mulByte_1_inst_00_o;
  wire [7:0] mulByte_2_inst_02_rhs;
  wire [7:0] mulByte_2_inst_02_o;
  wire [7:0] mulByte_2_inst_03_rhs;
  wire [7:0] mulByte_2_inst_03_o;
  wire [7:0] mulByte_2_inst_04_rhs;
  wire [7:0] mulByte_2_inst_04_o;
  wire [7:0] mulByte_0_inst_01_rhs;
  wire [7:0] mulByte_0_inst_01_o;
  wire [7:0] mulByte_1_inst_01_rhs;
  wire [7:0] mulByte_1_inst_01_o;
  wire [7:0] mulByte_1_inst_02_rhs;
  wire [7:0] mulByte_1_inst_02_o;
  wire [7:0] mulByte_2_inst_05_rhs;
  wire [7:0] mulByte_2_inst_05_o;
  wire [7:0] mulByte_2_inst_06_rhs;
  wire [7:0] mulByte_2_inst_06_o;
  wire [7:0] mulByte_0_inst_02_rhs;
  wire [7:0] mulByte_0_inst_02_o;
  wire [7:0] mulByte_0_inst_03_rhs;
  wire [7:0] mulByte_0_inst_03_o;
  wire [7:0] mulByte_1_inst_03_rhs;
  wire [7:0] mulByte_1_inst_03_o;
  wire [7:0] mulByte_2_inst_07_rhs;
  wire [7:0] mulByte_2_inst_07_o;
  wire [7:0] mulByte_2_inst_08_rhs;
  wire [7:0] mulByte_2_inst_08_o;
  wire [7:0] mulByte_2_inst_09_rhs;
  wire [7:0] mulByte_2_inst_09_o;
  wire [7:0] mulByte_0_inst_04_rhs;
  wire [7:0] mulByte_0_inst_04_o;
  wire [7:0] mulByte_1_inst_04_rhs;
  wire [7:0] mulByte_1_inst_04_o;
  wire [7:0] mulByte_2_inst_10_rhs;
  wire [7:0] mulByte_2_inst_10_o;
  wire [7:0] mulByte_2_inst_11_rhs;
  wire [7:0] mulByte_2_inst_11_o;
  wire [7:0] mulByte_2_inst_12_rhs;
  wire [7:0] mulByte_2_inst_12_o;
  wire [7:0] mulByte_0_inst_05_rhs;
  wire [7:0] mulByte_0_inst_05_o;
  wire [7:0] mulByte_1_inst_05_rhs;
  wire [7:0] mulByte_1_inst_05_o;
  wire [7:0] mulByte_1_inst_06_rhs;
  wire [7:0] mulByte_1_inst_06_o;
  wire [7:0] mulByte_2_inst_13_rhs;
  wire [7:0] mulByte_2_inst_13_o;
  wire [7:0] mulByte_2_inst_14_rhs;
  wire [7:0] mulByte_2_inst_14_o;
  wire [7:0] mulByte_0_inst_06_rhs;
  wire [7:0] mulByte_0_inst_06_o;
  wire [7:0] mulByte_0_inst_07_rhs;
  wire [7:0] mulByte_0_inst_07_o;
  wire [7:0] mulByte_1_inst_07_rhs;
  wire [7:0] mulByte_1_inst_07_o;
  wire [7:0] mulByte_2_inst_15_rhs;
  wire [7:0] mulByte_2_inst_15_o;
  wire [7:0] mulByte_2_inst_16_rhs;
  wire [7:0] mulByte_2_inst_16_o;
  wire [7:0] mulByte_2_inst_17_rhs;
  wire [7:0] mulByte_2_inst_17_o;
  wire [7:0] mulByte_0_inst_08_rhs;
  wire [7:0] mulByte_0_inst_08_o;
  wire [7:0] mulByte_1_inst_08_rhs;
  wire [7:0] mulByte_1_inst_08_o;
  wire [7:0] mulByte_2_inst_18_rhs;
  wire [7:0] mulByte_2_inst_18_o;
  wire [7:0] mulByte_2_inst_19_rhs;
  wire [7:0] mulByte_2_inst_19_o;
  wire [7:0] mulByte_2_inst_20_rhs;
  wire [7:0] mulByte_2_inst_20_o;
  wire [7:0] mulByte_0_inst_09_rhs;
  wire [7:0] mulByte_0_inst_09_o;
  wire [7:0] mulByte_1_inst_09_rhs;
  wire [7:0] mulByte_1_inst_09_o;
  wire [7:0] mulByte_1_inst_10_rhs;
  wire [7:0] mulByte_1_inst_10_o;
  wire [7:0] mulByte_2_inst_21_rhs;
  wire [7:0] mulByte_2_inst_21_o;
  wire [7:0] mulByte_2_inst_22_rhs;
  wire [7:0] mulByte_2_inst_22_o;
  wire [7:0] mulByte_0_inst_10_rhs;
  wire [7:0] mulByte_0_inst_10_o;
  wire [7:0] mulByte_0_inst_11_rhs;
  wire [7:0] mulByte_0_inst_11_o;
  wire [7:0] mulByte_1_inst_11_rhs;
  wire [7:0] mulByte_1_inst_11_o;
  wire [7:0] mulByte_2_inst_23_rhs;
  wire [7:0] mulByte_2_inst_23_o;
  wire [7:0] mulByte_2_inst_24_rhs;
  wire [7:0] mulByte_2_inst_24_o;
  wire [7:0] mulByte_2_inst_25_rhs;
  wire [7:0] mulByte_2_inst_25_o;
  wire [7:0] mulByte_0_inst_12_rhs;
  wire [7:0] mulByte_0_inst_12_o;
  wire [7:0] mulByte_1_inst_12_rhs;
  wire [7:0] mulByte_1_inst_12_o;
  wire [7:0] mulByte_2_inst_26_rhs;
  wire [7:0] mulByte_2_inst_26_o;
  wire [7:0] mulByte_2_inst_27_rhs;
  wire [7:0] mulByte_2_inst_27_o;
  wire [7:0] mulByte_2_inst_28_rhs;
  wire [7:0] mulByte_2_inst_28_o;
  wire [7:0] mulByte_0_inst_13_rhs;
  wire [7:0] mulByte_0_inst_13_o;
  wire [7:0] mulByte_1_inst_13_rhs;
  wire [7:0] mulByte_1_inst_13_o;
  wire [7:0] mulByte_1_inst_14_rhs;
  wire [7:0] mulByte_1_inst_14_o;
  wire [7:0] mulByte_2_inst_29_rhs;
  wire [7:0] mulByte_2_inst_29_o;
  wire [7:0] mulByte_2_inst_30_rhs;
  wire [7:0] mulByte_2_inst_30_o;
  wire [7:0] mulByte_0_inst_14_rhs;
  wire [7:0] mulByte_0_inst_14_o;
  mulByte_0 #(
    .lhs (8'h02)
  ) o_part_mulByte_0_inst(
    .rhs /*<--*/ (o_part_mulByte_0_inst_rhs),
    .o   /*-->*/ (o_part_mulByte_0_inst_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) o_part_mulByte_1_inst(
    .rhs /*<--*/ (o_part_mulByte_1_inst_rhs),
    .o   /*-->*/ (o_part_mulByte_1_inst_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) o_part_mulByte_2_inst(
    .rhs /*<--*/ (o_part_mulByte_2_inst_rhs),
    .o   /*-->*/ (o_part_mulByte_2_inst_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_00(
    .rhs /*<--*/ (mulByte_2_inst_00_rhs),
    .o   /*-->*/ (mulByte_2_inst_00_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_01(
    .rhs /*<--*/ (mulByte_2_inst_01_rhs),
    .o   /*-->*/ (mulByte_2_inst_01_o)
  );
  mulByte_0 #(
    .lhs (8'h02)
  ) mulByte_0_inst_00(
    .rhs /*<--*/ (mulByte_0_inst_00_rhs),
    .o   /*-->*/ (mulByte_0_inst_00_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) mulByte_1_inst_00(
    .rhs /*<--*/ (mulByte_1_inst_00_rhs),
    .o   /*-->*/ (mulByte_1_inst_00_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_02(
    .rhs /*<--*/ (mulByte_2_inst_02_rhs),
    .o   /*-->*/ (mulByte_2_inst_02_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_03(
    .rhs /*<--*/ (mulByte_2_inst_03_rhs),
    .o   /*-->*/ (mulByte_2_inst_03_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_04(
    .rhs /*<--*/ (mulByte_2_inst_04_rhs),
    .o   /*-->*/ (mulByte_2_inst_04_o)
  );
  mulByte_0 #(
    .lhs (8'h02)
  ) mulByte_0_inst_01(
    .rhs /*<--*/ (mulByte_0_inst_01_rhs),
    .o   /*-->*/ (mulByte_0_inst_01_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) mulByte_1_inst_01(
    .rhs /*<--*/ (mulByte_1_inst_01_rhs),
    .o   /*-->*/ (mulByte_1_inst_01_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) mulByte_1_inst_02(
    .rhs /*<--*/ (mulByte_1_inst_02_rhs),
    .o   /*-->*/ (mulByte_1_inst_02_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_05(
    .rhs /*<--*/ (mulByte_2_inst_05_rhs),
    .o   /*-->*/ (mulByte_2_inst_05_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_06(
    .rhs /*<--*/ (mulByte_2_inst_06_rhs),
    .o   /*-->*/ (mulByte_2_inst_06_o)
  );
  mulByte_0 #(
    .lhs (8'h02)
  ) mulByte_0_inst_02(
    .rhs /*<--*/ (mulByte_0_inst_02_rhs),
    .o   /*-->*/ (mulByte_0_inst_02_o)
  );
  mulByte_0 #(
    .lhs (8'h02)
  ) mulByte_0_inst_03(
    .rhs /*<--*/ (mulByte_0_inst_03_rhs),
    .o   /*-->*/ (mulByte_0_inst_03_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) mulByte_1_inst_03(
    .rhs /*<--*/ (mulByte_1_inst_03_rhs),
    .o   /*-->*/ (mulByte_1_inst_03_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_07(
    .rhs /*<--*/ (mulByte_2_inst_07_rhs),
    .o   /*-->*/ (mulByte_2_inst_07_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_08(
    .rhs /*<--*/ (mulByte_2_inst_08_rhs),
    .o   /*-->*/ (mulByte_2_inst_08_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_09(
    .rhs /*<--*/ (mulByte_2_inst_09_rhs),
    .o   /*-->*/ (mulByte_2_inst_09_o)
  );
  mulByte_0 #(
    .lhs (8'h02)
  ) mulByte_0_inst_04(
    .rhs /*<--*/ (mulByte_0_inst_04_rhs),
    .o   /*-->*/ (mulByte_0_inst_04_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) mulByte_1_inst_04(
    .rhs /*<--*/ (mulByte_1_inst_04_rhs),
    .o   /*-->*/ (mulByte_1_inst_04_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_10(
    .rhs /*<--*/ (mulByte_2_inst_10_rhs),
    .o   /*-->*/ (mulByte_2_inst_10_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_11(
    .rhs /*<--*/ (mulByte_2_inst_11_rhs),
    .o   /*-->*/ (mulByte_2_inst_11_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_12(
    .rhs /*<--*/ (mulByte_2_inst_12_rhs),
    .o   /*-->*/ (mulByte_2_inst_12_o)
  );
  mulByte_0 #(
    .lhs (8'h02)
  ) mulByte_0_inst_05(
    .rhs /*<--*/ (mulByte_0_inst_05_rhs),
    .o   /*-->*/ (mulByte_0_inst_05_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) mulByte_1_inst_05(
    .rhs /*<--*/ (mulByte_1_inst_05_rhs),
    .o   /*-->*/ (mulByte_1_inst_05_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) mulByte_1_inst_06(
    .rhs /*<--*/ (mulByte_1_inst_06_rhs),
    .o   /*-->*/ (mulByte_1_inst_06_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_13(
    .rhs /*<--*/ (mulByte_2_inst_13_rhs),
    .o   /*-->*/ (mulByte_2_inst_13_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_14(
    .rhs /*<--*/ (mulByte_2_inst_14_rhs),
    .o   /*-->*/ (mulByte_2_inst_14_o)
  );
  mulByte_0 #(
    .lhs (8'h02)
  ) mulByte_0_inst_06(
    .rhs /*<--*/ (mulByte_0_inst_06_rhs),
    .o   /*-->*/ (mulByte_0_inst_06_o)
  );
  mulByte_0 #(
    .lhs (8'h02)
  ) mulByte_0_inst_07(
    .rhs /*<--*/ (mulByte_0_inst_07_rhs),
    .o   /*-->*/ (mulByte_0_inst_07_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) mulByte_1_inst_07(
    .rhs /*<--*/ (mulByte_1_inst_07_rhs),
    .o   /*-->*/ (mulByte_1_inst_07_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_15(
    .rhs /*<--*/ (mulByte_2_inst_15_rhs),
    .o   /*-->*/ (mulByte_2_inst_15_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_16(
    .rhs /*<--*/ (mulByte_2_inst_16_rhs),
    .o   /*-->*/ (mulByte_2_inst_16_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_17(
    .rhs /*<--*/ (mulByte_2_inst_17_rhs),
    .o   /*-->*/ (mulByte_2_inst_17_o)
  );
  mulByte_0 #(
    .lhs (8'h02)
  ) mulByte_0_inst_08(
    .rhs /*<--*/ (mulByte_0_inst_08_rhs),
    .o   /*-->*/ (mulByte_0_inst_08_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) mulByte_1_inst_08(
    .rhs /*<--*/ (mulByte_1_inst_08_rhs),
    .o   /*-->*/ (mulByte_1_inst_08_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_18(
    .rhs /*<--*/ (mulByte_2_inst_18_rhs),
    .o   /*-->*/ (mulByte_2_inst_18_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_19(
    .rhs /*<--*/ (mulByte_2_inst_19_rhs),
    .o   /*-->*/ (mulByte_2_inst_19_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_20(
    .rhs /*<--*/ (mulByte_2_inst_20_rhs),
    .o   /*-->*/ (mulByte_2_inst_20_o)
  );
  mulByte_0 #(
    .lhs (8'h02)
  ) mulByte_0_inst_09(
    .rhs /*<--*/ (mulByte_0_inst_09_rhs),
    .o   /*-->*/ (mulByte_0_inst_09_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) mulByte_1_inst_09(
    .rhs /*<--*/ (mulByte_1_inst_09_rhs),
    .o   /*-->*/ (mulByte_1_inst_09_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) mulByte_1_inst_10(
    .rhs /*<--*/ (mulByte_1_inst_10_rhs),
    .o   /*-->*/ (mulByte_1_inst_10_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_21(
    .rhs /*<--*/ (mulByte_2_inst_21_rhs),
    .o   /*-->*/ (mulByte_2_inst_21_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_22(
    .rhs /*<--*/ (mulByte_2_inst_22_rhs),
    .o   /*-->*/ (mulByte_2_inst_22_o)
  );
  mulByte_0 #(
    .lhs (8'h02)
  ) mulByte_0_inst_10(
    .rhs /*<--*/ (mulByte_0_inst_10_rhs),
    .o   /*-->*/ (mulByte_0_inst_10_o)
  );
  mulByte_0 #(
    .lhs (8'h02)
  ) mulByte_0_inst_11(
    .rhs /*<--*/ (mulByte_0_inst_11_rhs),
    .o   /*-->*/ (mulByte_0_inst_11_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) mulByte_1_inst_11(
    .rhs /*<--*/ (mulByte_1_inst_11_rhs),
    .o   /*-->*/ (mulByte_1_inst_11_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_23(
    .rhs /*<--*/ (mulByte_2_inst_23_rhs),
    .o   /*-->*/ (mulByte_2_inst_23_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_24(
    .rhs /*<--*/ (mulByte_2_inst_24_rhs),
    .o   /*-->*/ (mulByte_2_inst_24_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_25(
    .rhs /*<--*/ (mulByte_2_inst_25_rhs),
    .o   /*-->*/ (mulByte_2_inst_25_o)
  );
  mulByte_0 #(
    .lhs (8'h02)
  ) mulByte_0_inst_12(
    .rhs /*<--*/ (mulByte_0_inst_12_rhs),
    .o   /*-->*/ (mulByte_0_inst_12_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) mulByte_1_inst_12(
    .rhs /*<--*/ (mulByte_1_inst_12_rhs),
    .o   /*-->*/ (mulByte_1_inst_12_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_26(
    .rhs /*<--*/ (mulByte_2_inst_26_rhs),
    .o   /*-->*/ (mulByte_2_inst_26_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_27(
    .rhs /*<--*/ (mulByte_2_inst_27_rhs),
    .o   /*-->*/ (mulByte_2_inst_27_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_28(
    .rhs /*<--*/ (mulByte_2_inst_28_rhs),
    .o   /*-->*/ (mulByte_2_inst_28_o)
  );
  mulByte_0 #(
    .lhs (8'h02)
  ) mulByte_0_inst_13(
    .rhs /*<--*/ (mulByte_0_inst_13_rhs),
    .o   /*-->*/ (mulByte_0_inst_13_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) mulByte_1_inst_13(
    .rhs /*<--*/ (mulByte_1_inst_13_rhs),
    .o   /*-->*/ (mulByte_1_inst_13_o)
  );
  mulByte_1 #(
    .lhs (8'h03)
  ) mulByte_1_inst_14(
    .rhs /*<--*/ (mulByte_1_inst_14_rhs),
    .o   /*-->*/ (mulByte_1_inst_14_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_29(
    .rhs /*<--*/ (mulByte_2_inst_29_rhs),
    .o   /*-->*/ (mulByte_2_inst_29_o)
  );
  mulByte_2 #(
    .lhs (8'h01)
  ) mulByte_2_inst_30(
    .rhs /*<--*/ (mulByte_2_inst_30_rhs),
    .o   /*-->*/ (mulByte_2_inst_30_o)
  );
  mulByte_0 #(
    .lhs (8'h02)
  ) mulByte_0_inst_14(
    .rhs /*<--*/ (mulByte_0_inst_14_rhs),
    .o   /*-->*/ (mulByte_0_inst_14_o)
  );
  assign o_part_mulByte_0_inst_rhs = state[0][0];
  assign o_part_mulByte_1_inst_rhs = state[0][1];
  assign o_part_mulByte_2_inst_rhs = state[0][2];
  assign mulByte_2_inst_00_rhs = state[0][3];
  assign mulByte_2_inst_01_rhs = state[0][0];
  assign mulByte_0_inst_00_rhs = state[0][1];
  assign mulByte_1_inst_00_rhs = state[0][2];
  assign mulByte_2_inst_02_rhs = state[0][3];
  assign mulByte_2_inst_03_rhs = state[0][0];
  assign mulByte_2_inst_04_rhs = state[0][1];
  assign mulByte_0_inst_01_rhs = state[0][2];
  assign mulByte_1_inst_01_rhs = state[0][3];
  assign mulByte_1_inst_02_rhs = state[0][0];
  assign mulByte_2_inst_05_rhs = state[0][1];
  assign mulByte_2_inst_06_rhs = state[0][2];
  assign mulByte_0_inst_02_rhs = state[0][3];
  assign mulByte_0_inst_03_rhs = state[1][0];
  assign mulByte_1_inst_03_rhs = state[1][1];
  assign mulByte_2_inst_07_rhs = state[1][2];
  assign mulByte_2_inst_08_rhs = state[1][3];
  assign mulByte_2_inst_09_rhs = state[1][0];
  assign mulByte_0_inst_04_rhs = state[1][1];
  assign mulByte_1_inst_04_rhs = state[1][2];
  assign mulByte_2_inst_10_rhs = state[1][3];
  assign mulByte_2_inst_11_rhs = state[1][0];
  assign mulByte_2_inst_12_rhs = state[1][1];
  assign mulByte_0_inst_05_rhs = state[1][2];
  assign mulByte_1_inst_05_rhs = state[1][3];
  assign mulByte_1_inst_06_rhs = state[1][0];
  assign mulByte_2_inst_13_rhs = state[1][1];
  assign mulByte_2_inst_14_rhs = state[1][2];
  assign mulByte_0_inst_06_rhs = state[1][3];
  assign mulByte_0_inst_07_rhs = state[2][0];
  assign mulByte_1_inst_07_rhs = state[2][1];
  assign mulByte_2_inst_15_rhs = state[2][2];
  assign mulByte_2_inst_16_rhs = state[2][3];
  assign mulByte_2_inst_17_rhs = state[2][0];
  assign mulByte_0_inst_08_rhs = state[2][1];
  assign mulByte_1_inst_08_rhs = state[2][2];
  assign mulByte_2_inst_18_rhs = state[2][3];
  assign mulByte_2_inst_19_rhs = state[2][0];
  assign mulByte_2_inst_20_rhs = state[2][1];
  assign mulByte_0_inst_09_rhs = state[2][2];
  assign mulByte_1_inst_09_rhs = state[2][3];
  assign mulByte_1_inst_10_rhs = state[2][0];
  assign mulByte_2_inst_21_rhs = state[2][1];
  assign mulByte_2_inst_22_rhs = state[2][2];
  assign mulByte_0_inst_10_rhs = state[2][3];
  assign mulByte_0_inst_11_rhs = state[3][0];
  assign mulByte_1_inst_11_rhs = state[3][1];
  assign mulByte_2_inst_23_rhs = state[3][2];
  assign mulByte_2_inst_24_rhs = state[3][3];
  assign mulByte_2_inst_25_rhs = state[3][0];
  assign mulByte_0_inst_12_rhs = state[3][1];
  assign mulByte_1_inst_12_rhs = state[3][2];
  assign mulByte_2_inst_26_rhs = state[3][3];
  assign mulByte_2_inst_27_rhs = state[3][0];
  assign mulByte_2_inst_28_rhs = state[3][1];
  assign mulByte_0_inst_13_rhs = state[3][2];
  assign mulByte_1_inst_13_rhs = state[3][3];
  assign mulByte_1_inst_14_rhs = state[3][0];
  assign mulByte_2_inst_29_rhs = state[3][1];
  assign mulByte_2_inst_30_rhs = state[3][2];
  assign mulByte_0_inst_14_rhs = state[3][3];
  assign o = '{
    '{
      ((o_part_mulByte_0_inst_o ^ o_part_mulByte_1_inst_o) ^ o_part_mulByte_2_inst_o) ^ mulByte_2_inst_00_o,
      ((mulByte_2_inst_01_o ^ mulByte_0_inst_00_o) ^ mulByte_1_inst_00_o) ^ mulByte_2_inst_02_o,
      ((mulByte_2_inst_03_o ^ mulByte_2_inst_04_o) ^ mulByte_0_inst_01_o) ^ mulByte_1_inst_01_o,
      ((mulByte_1_inst_02_o ^ mulByte_2_inst_05_o) ^ mulByte_2_inst_06_o) ^ mulByte_0_inst_02_o
    },
    '{
      ((mulByte_0_inst_03_o ^ mulByte_1_inst_03_o) ^ mulByte_2_inst_07_o) ^ mulByte_2_inst_08_o,
      ((mulByte_2_inst_09_o ^ mulByte_0_inst_04_o) ^ mulByte_1_inst_04_o) ^ mulByte_2_inst_10_o,
      ((mulByte_2_inst_11_o ^ mulByte_2_inst_12_o) ^ mulByte_0_inst_05_o) ^ mulByte_1_inst_05_o,
      ((mulByte_1_inst_06_o ^ mulByte_2_inst_13_o) ^ mulByte_2_inst_14_o) ^ mulByte_0_inst_06_o
    },
    '{
      ((mulByte_0_inst_07_o ^ mulByte_1_inst_07_o) ^ mulByte_2_inst_15_o) ^ mulByte_2_inst_16_o,
      ((mulByte_2_inst_17_o ^ mulByte_0_inst_08_o) ^ mulByte_1_inst_08_o) ^ mulByte_2_inst_18_o,
      ((mulByte_2_inst_19_o ^ mulByte_2_inst_20_o) ^ mulByte_0_inst_09_o) ^ mulByte_1_inst_09_o,
      ((mulByte_1_inst_10_o ^ mulByte_2_inst_21_o) ^ mulByte_2_inst_22_o) ^ mulByte_0_inst_10_o
    },
    '{
      ((mulByte_0_inst_11_o ^ mulByte_1_inst_11_o) ^ mulByte_2_inst_23_o) ^ mulByte_2_inst_24_o,
      ((mulByte_2_inst_25_o ^ mulByte_0_inst_12_o) ^ mulByte_1_inst_12_o) ^ mulByte_2_inst_26_o,
      ((mulByte_2_inst_27_o ^ mulByte_2_inst_28_o) ^ mulByte_0_inst_13_o) ^ mulByte_1_inst_13_o,
      ((mulByte_1_inst_14_o ^ mulByte_2_inst_29_o) ^ mulByte_2_inst_30_o) ^ mulByte_0_inst_14_o
    }
  };
endmodule
