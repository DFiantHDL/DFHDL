`ifndef UART_TX_DEFS
`define UART_TX_DEFS

`endif
`ifndef UART_TX_DEFS_MODULE
`define UART_TX_DEFS_MODULE
`else

`undef UART_TX_DEFS_MODULE
`endif

