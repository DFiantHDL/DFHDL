`ifndef ALU_DEFS
`define ALU_DEFS
`define ALUSel_ADD 0
`define ALUSel_SUB 1
`define ALUSel_SLL 2
`define ALUSel_SRL 3
`define ALUSel_SRA 4
`define ALUSel_AND 5
`define ALUSel_OR 6
`define ALUSel_XOR 7
`define ALUSel_SLT 8
`define ALUSel_SLTU 9
`define ALUSel_COPY1 10

`endif
