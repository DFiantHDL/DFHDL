`ifndef FULLADDERN_DEFS
`define FULLADDERN_DEFS
`endif
