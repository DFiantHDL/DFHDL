`ifndef LRSHIFTDIRECT_DEFS
`define LRSHIFTDIRECT_DEFS
`define ShiftDir_Left 0
`define ShiftDir_Right 1

`endif
