`ifndef LRSHIFTDIRECT_DEFS
`define LRSHIFTDIRECT_DEFS
typedef enum logic [0:0] {
  ShiftDir_Left  = 0,
  ShiftDir_Right = 1
} t_enum_ShiftDir;
`endif
