`ifndef REGFILE_DEFS
`define REGFILE_DEFS

`endif
