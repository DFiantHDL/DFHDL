`ifndef FULLADDER1_DEFS
`define FULLADDER1_DEFS

`endif
`ifndef FULLADDER1_DEFS_MODULE
`define FULLADDER1_DEFS_MODULE
`else

`undef FULLADDER1_DEFS_MODULE
`endif

