`ifndef LEFTSHIFTGEN_DEFS
`define LEFTSHIFTGEN_DEFS

`endif
