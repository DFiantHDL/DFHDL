`ifndef CIPHER_DEFS
`define CIPHER_DEFS
typedef logic [7:0] t_opaque_AESByte;
typedef t_opaque_AESByte t_opaque_AESWord [0:3];
typedef t_opaque_AESWord t_opaque_AESKey [0:3];
typedef t_opaque_AESWord t_opaque_AESData [0:3];
typedef t_opaque_AESWord t_opaque_AESKeySchedule [0:43];
typedef t_opaque_AESWord t_opaque_AESState [0:3];
typedef t_opaque_AESWord t_opaque_AESRoundKey [0:3];
parameter logic [7:0] sboxLookupTable [0:255] = '{
    0: 8'h63,   1: 8'h7c,   2: 8'h77,   3: 8'h7b,   4: 8'hf2,   5: 8'h6b,   6: 8'h6f,   7: 8'hc5,
    8: 8'h30,   9: 8'h01,  10: 8'h67,  11: 8'h2b,  12: 8'hfe,  13: 8'hd7,  14: 8'hab,  15: 8'h76,
   16: 8'hca,  17: 8'h82,  18: 8'hc9,  19: 8'h7d,  20: 8'hfa,  21: 8'h59,  22: 8'h47,  23: 8'hf0,
   24: 8'had,  25: 8'hd4,  26: 8'ha2,  27: 8'haf,  28: 8'h9c,  29: 8'ha4,  30: 8'h72,  31: 8'hc0,
   32: 8'hb7,  33: 8'hfd,  34: 8'h93,  35: 8'h26,  36: 8'h36,  37: 8'h3f,  38: 8'hf7,  39: 8'hcc,
   40: 8'h34,  41: 8'ha5,  42: 8'he5,  43: 8'hf1,  44: 8'h71,  45: 8'hd8,  46: 8'h31,  47: 8'h15,
   48: 8'h04,  49: 8'hc7,  50: 8'h23,  51: 8'hc3,  52: 8'h18,  53: 8'h96,  54: 8'h05,  55: 8'h9a,
   56: 8'h07,  57: 8'h12,  58: 8'h80,  59: 8'he2,  60: 8'heb,  61: 8'h27,  62: 8'hb2,  63: 8'h75,
   64: 8'h09,  65: 8'h83,  66: 8'h2c,  67: 8'h1a,  68: 8'h1b,  69: 8'h6e,  70: 8'h5a,  71: 8'ha0,
   72: 8'h52,  73: 8'h3b,  74: 8'hd6,  75: 8'hb3,  76: 8'h29,  77: 8'he3,  78: 8'h2f,  79: 8'h84,
   80: 8'h53,  81: 8'hd1,  82: 8'h00,  83: 8'hed,  84: 8'h20,  85: 8'hfc,  86: 8'hb1,  87: 8'h5b,
   88: 8'h6a,  89: 8'hcb,  90: 8'hbe,  91: 8'h39,  92: 8'h4a,  93: 8'h4c,  94: 8'h58,  95: 8'hcf,
   96: 8'hd0,  97: 8'hef,  98: 8'haa,  99: 8'hfb, 100: 8'h43, 101: 8'h4d, 102: 8'h33, 103: 8'h85,
  104: 8'h45, 105: 8'hf9, 106: 8'h02, 107: 8'h7f, 108: 8'h50, 109: 8'h3c, 110: 8'h9f, 111: 8'ha8,
  112: 8'h51, 113: 8'ha3, 114: 8'h40, 115: 8'h8f, 116: 8'h92, 117: 8'h9d, 118: 8'h38, 119: 8'hf5,
  120: 8'hbc, 121: 8'hb6, 122: 8'hda, 123: 8'h21, 124: 8'h10, 125: 8'hff, 126: 8'hf3, 127: 8'hd2,
  128: 8'hcd, 129: 8'h0c, 130: 8'h13, 131: 8'hec, 132: 8'h5f, 133: 8'h97, 134: 8'h44, 135: 8'h17,
  136: 8'hc4, 137: 8'ha7, 138: 8'h7e, 139: 8'h3d, 140: 8'h64, 141: 8'h5d, 142: 8'h19, 143: 8'h73,
  144: 8'h60, 145: 8'h81, 146: 8'h4f, 147: 8'hdc, 148: 8'h22, 149: 8'h2a, 150: 8'h90, 151: 8'h88,
  152: 8'h46, 153: 8'hee, 154: 8'hb8, 155: 8'h14, 156: 8'hde, 157: 8'h5e, 158: 8'h0b, 159: 8'hdb,
  160: 8'he0, 161: 8'h32, 162: 8'h3a, 163: 8'h0a, 164: 8'h49, 165: 8'h06, 166: 8'h24, 167: 8'h5c,
  168: 8'hc2, 169: 8'hd3, 170: 8'hac, 171: 8'h62, 172: 8'h91, 173: 8'h95, 174: 8'he4, 175: 8'h79,
  176: 8'he7, 177: 8'hc8, 178: 8'h37, 179: 8'h6d, 180: 8'h8d, 181: 8'hd5, 182: 8'h4e, 183: 8'ha9,
  184: 8'h6c, 185: 8'h56, 186: 8'hf4, 187: 8'hea, 188: 8'h65, 189: 8'h7a, 190: 8'hae, 191: 8'h08,
  192: 8'hba, 193: 8'h78, 194: 8'h25, 195: 8'h2e, 196: 8'h1c, 197: 8'ha6, 198: 8'hb4, 199: 8'hc6,
  200: 8'he8, 201: 8'hdd, 202: 8'h74, 203: 8'h1f, 204: 8'h4b, 205: 8'hbd, 206: 8'h8b, 207: 8'h8a,
  208: 8'h70, 209: 8'h3e, 210: 8'hb5, 211: 8'h66, 212: 8'h48, 213: 8'h03, 214: 8'hf6, 215: 8'h0e,
  216: 8'h61, 217: 8'h35, 218: 8'h57, 219: 8'hb9, 220: 8'h86, 221: 8'hc1, 222: 8'h1d, 223: 8'h9e,
  224: 8'he1, 225: 8'hf8, 226: 8'h98, 227: 8'h11, 228: 8'h69, 229: 8'hd9, 230: 8'h8e, 231: 8'h94,
  232: 8'h9b, 233: 8'h1e, 234: 8'h87, 235: 8'he9, 236: 8'hce, 237: 8'h55, 238: 8'h28, 239: 8'hdf,
  240: 8'h8c, 241: 8'ha1, 242: 8'h89, 243: 8'h0d, 244: 8'hbf, 245: 8'he6, 246: 8'h42, 247: 8'h68,
  248: 8'h41, 249: 8'h99, 250: 8'h2d, 251: 8'h0f, 252: 8'hb0, 253: 8'h54, 254: 8'hbb, 255: 8'h16
};
parameter t_opaque_AESWord Rcon [0:10] = '{
   0: '{0: 8'h00, 1: 8'h00, 2: 8'h00, 3: 8'h00},
   1: '{0: 8'h01, 1: 8'h00, 2: 8'h00, 3: 8'h00},
   2: '{0: 8'h02, 1: 8'h00, 2: 8'h00, 3: 8'h00},
   3: '{0: 8'h04, 1: 8'h00, 2: 8'h00, 3: 8'h00},
   4: '{0: 8'h08, 1: 8'h00, 2: 8'h00, 3: 8'h00},
   5: '{0: 8'h10, 1: 8'h00, 2: 8'h00, 3: 8'h00},
   6: '{0: 8'h20, 1: 8'h00, 2: 8'h00, 3: 8'h00},
   7: '{0: 8'h40, 1: 8'h00, 2: 8'h00, 3: 8'h00},
   8: '{0: 8'h80, 1: 8'h00, 2: 8'h00, 3: 8'h00},
   9: '{0: 8'h1b, 1: 8'h00, 2: 8'h00, 3: 8'h00},
  10: '{0: 8'h36, 1: 8'h00, 2: 8'h00, 3: 8'h00}
};
`endif
