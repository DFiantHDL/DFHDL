`ifndef LEFTSHIFTBASIC_DEFS
`define LEFTSHIFTBASIC_DEFS

`endif
