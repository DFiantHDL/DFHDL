library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.dfhdl_pkg.all;

package TrueDPR_pkg is
end package TrueDPR_pkg;

package body TrueDPR_pkg is
end package body TrueDPR_pkg;
