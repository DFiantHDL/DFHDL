`ifndef LEFTSHIFTBASIC_DEFS
`define LEFTSHIFTBASIC_DEFS

`endif
`ifndef LEFTSHIFTBASIC_DEFS_MODULE
`define LEFTSHIFTBASIC_DEFS_MODULE
`else

`undef LEFTSHIFTBASIC_DEFS_MODULE
`endif

