library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.dfhdl_pkg.all;

package Counter_pkg is

end package Counter_pkg;

package body Counter_pkg is

end package body Counter_pkg;
