library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.dfhdl_pkg.all;

package UART_Tx_pkg is

end package UART_Tx_pkg;

package body UART_Tx_pkg is

end package body UART_Tx_pkg;
