`ifndef FULLADDER1_DEFS
`define FULLADDER1_DEFS

`endif
