library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.dfhdl_pkg.all;

package FullAdder1_pkg is

end package FullAdder1_pkg;

package body FullAdder1_pkg is

end package body FullAdder1_pkg;
