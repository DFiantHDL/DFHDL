`ifndef LEFTSHIFT2_DEFS
`define LEFTSHIFT2_DEFS

`endif
