`ifndef UART_TX_DEFS
`define UART_TX_DEFS

`endif
