`ifndef REGFILE_DEFS
`define REGFILE_DEFS
`endif
`ifndef REGFILE_DEFS_MODULE
`define REGFILE_DEFS_MODULE
`else
`undef REGFILE_DEFS_MODULE
`endif
