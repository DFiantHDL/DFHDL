library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.dfhdl_pkg.all;
use work.CipherNoOpaques_pkg.all;

entity mixColumns is
port (
  state : in  t_opaque_AESState;
  o     : out t_opaque_AESState
);
end mixColumns;

architecture mixColumns_arch of mixColumns is
  signal o_part_mulByte_0_inst_rhs : t_opaque_AESByte;
  signal o_part_mulByte_0_inst_o   : t_opaque_AESByte;
  signal o_part_mulByte_1_inst_rhs : t_opaque_AESByte;
  signal o_part_mulByte_1_inst_o   : t_opaque_AESByte;
  signal o_part_mulByte_2_inst_rhs : t_opaque_AESByte;
  signal o_part_mulByte_2_inst_o   : t_opaque_AESByte;
  signal mulByte_2_inst_00_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_00_o       : t_opaque_AESByte;
  signal mulByte_2_inst_01_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_01_o       : t_opaque_AESByte;
  signal mulByte_0_inst_00_rhs     : t_opaque_AESByte;
  signal mulByte_0_inst_00_o       : t_opaque_AESByte;
  signal mulByte_1_inst_00_rhs     : t_opaque_AESByte;
  signal mulByte_1_inst_00_o       : t_opaque_AESByte;
  signal mulByte_2_inst_02_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_02_o       : t_opaque_AESByte;
  signal mulByte_2_inst_03_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_03_o       : t_opaque_AESByte;
  signal mulByte_2_inst_04_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_04_o       : t_opaque_AESByte;
  signal mulByte_0_inst_01_rhs     : t_opaque_AESByte;
  signal mulByte_0_inst_01_o       : t_opaque_AESByte;
  signal mulByte_1_inst_01_rhs     : t_opaque_AESByte;
  signal mulByte_1_inst_01_o       : t_opaque_AESByte;
  signal mulByte_1_inst_02_rhs     : t_opaque_AESByte;
  signal mulByte_1_inst_02_o       : t_opaque_AESByte;
  signal mulByte_2_inst_05_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_05_o       : t_opaque_AESByte;
  signal mulByte_2_inst_06_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_06_o       : t_opaque_AESByte;
  signal mulByte_0_inst_02_rhs     : t_opaque_AESByte;
  signal mulByte_0_inst_02_o       : t_opaque_AESByte;
  signal mulByte_0_inst_03_rhs     : t_opaque_AESByte;
  signal mulByte_0_inst_03_o       : t_opaque_AESByte;
  signal mulByte_1_inst_03_rhs     : t_opaque_AESByte;
  signal mulByte_1_inst_03_o       : t_opaque_AESByte;
  signal mulByte_2_inst_07_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_07_o       : t_opaque_AESByte;
  signal mulByte_2_inst_08_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_08_o       : t_opaque_AESByte;
  signal mulByte_2_inst_09_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_09_o       : t_opaque_AESByte;
  signal mulByte_0_inst_04_rhs     : t_opaque_AESByte;
  signal mulByte_0_inst_04_o       : t_opaque_AESByte;
  signal mulByte_1_inst_04_rhs     : t_opaque_AESByte;
  signal mulByte_1_inst_04_o       : t_opaque_AESByte;
  signal mulByte_2_inst_10_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_10_o       : t_opaque_AESByte;
  signal mulByte_2_inst_11_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_11_o       : t_opaque_AESByte;
  signal mulByte_2_inst_12_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_12_o       : t_opaque_AESByte;
  signal mulByte_0_inst_05_rhs     : t_opaque_AESByte;
  signal mulByte_0_inst_05_o       : t_opaque_AESByte;
  signal mulByte_1_inst_05_rhs     : t_opaque_AESByte;
  signal mulByte_1_inst_05_o       : t_opaque_AESByte;
  signal mulByte_1_inst_06_rhs     : t_opaque_AESByte;
  signal mulByte_1_inst_06_o       : t_opaque_AESByte;
  signal mulByte_2_inst_13_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_13_o       : t_opaque_AESByte;
  signal mulByte_2_inst_14_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_14_o       : t_opaque_AESByte;
  signal mulByte_0_inst_06_rhs     : t_opaque_AESByte;
  signal mulByte_0_inst_06_o       : t_opaque_AESByte;
  signal mulByte_0_inst_07_rhs     : t_opaque_AESByte;
  signal mulByte_0_inst_07_o       : t_opaque_AESByte;
  signal mulByte_1_inst_07_rhs     : t_opaque_AESByte;
  signal mulByte_1_inst_07_o       : t_opaque_AESByte;
  signal mulByte_2_inst_15_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_15_o       : t_opaque_AESByte;
  signal mulByte_2_inst_16_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_16_o       : t_opaque_AESByte;
  signal mulByte_2_inst_17_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_17_o       : t_opaque_AESByte;
  signal mulByte_0_inst_08_rhs     : t_opaque_AESByte;
  signal mulByte_0_inst_08_o       : t_opaque_AESByte;
  signal mulByte_1_inst_08_rhs     : t_opaque_AESByte;
  signal mulByte_1_inst_08_o       : t_opaque_AESByte;
  signal mulByte_2_inst_18_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_18_o       : t_opaque_AESByte;
  signal mulByte_2_inst_19_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_19_o       : t_opaque_AESByte;
  signal mulByte_2_inst_20_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_20_o       : t_opaque_AESByte;
  signal mulByte_0_inst_09_rhs     : t_opaque_AESByte;
  signal mulByte_0_inst_09_o       : t_opaque_AESByte;
  signal mulByte_1_inst_09_rhs     : t_opaque_AESByte;
  signal mulByte_1_inst_09_o       : t_opaque_AESByte;
  signal mulByte_1_inst_10_rhs     : t_opaque_AESByte;
  signal mulByte_1_inst_10_o       : t_opaque_AESByte;
  signal mulByte_2_inst_21_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_21_o       : t_opaque_AESByte;
  signal mulByte_2_inst_22_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_22_o       : t_opaque_AESByte;
  signal mulByte_0_inst_10_rhs     : t_opaque_AESByte;
  signal mulByte_0_inst_10_o       : t_opaque_AESByte;
  signal mulByte_0_inst_11_rhs     : t_opaque_AESByte;
  signal mulByte_0_inst_11_o       : t_opaque_AESByte;
  signal mulByte_1_inst_11_rhs     : t_opaque_AESByte;
  signal mulByte_1_inst_11_o       : t_opaque_AESByte;
  signal mulByte_2_inst_23_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_23_o       : t_opaque_AESByte;
  signal mulByte_2_inst_24_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_24_o       : t_opaque_AESByte;
  signal mulByte_2_inst_25_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_25_o       : t_opaque_AESByte;
  signal mulByte_0_inst_12_rhs     : t_opaque_AESByte;
  signal mulByte_0_inst_12_o       : t_opaque_AESByte;
  signal mulByte_1_inst_12_rhs     : t_opaque_AESByte;
  signal mulByte_1_inst_12_o       : t_opaque_AESByte;
  signal mulByte_2_inst_26_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_26_o       : t_opaque_AESByte;
  signal mulByte_2_inst_27_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_27_o       : t_opaque_AESByte;
  signal mulByte_2_inst_28_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_28_o       : t_opaque_AESByte;
  signal mulByte_0_inst_13_rhs     : t_opaque_AESByte;
  signal mulByte_0_inst_13_o       : t_opaque_AESByte;
  signal mulByte_1_inst_13_rhs     : t_opaque_AESByte;
  signal mulByte_1_inst_13_o       : t_opaque_AESByte;
  signal mulByte_1_inst_14_rhs     : t_opaque_AESByte;
  signal mulByte_1_inst_14_o       : t_opaque_AESByte;
  signal mulByte_2_inst_29_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_29_o       : t_opaque_AESByte;
  signal mulByte_2_inst_30_rhs     : t_opaque_AESByte;
  signal mulByte_2_inst_30_o       : t_opaque_AESByte;
  signal mulByte_0_inst_14_rhs     : t_opaque_AESByte;
  signal mulByte_0_inst_14_o       : t_opaque_AESByte;
begin
  o_part_mulByte_0_inst : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => o_part_mulByte_0_inst_rhs,
    o   => o_part_mulByte_0_inst_o
  );
  o_part_mulByte_1_inst : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => o_part_mulByte_1_inst_rhs,
    o   => o_part_mulByte_1_inst_o
  );
  o_part_mulByte_2_inst : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => o_part_mulByte_2_inst_rhs,
    o   => o_part_mulByte_2_inst_o
  );
  mulByte_2_inst_00 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_00_rhs,
    o   => mulByte_2_inst_00_o
  );
  mulByte_2_inst_01 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_01_rhs,
    o   => mulByte_2_inst_01_o
  );
  mulByte_0_inst_00 : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => mulByte_0_inst_00_rhs,
    o   => mulByte_0_inst_00_o
  );
  mulByte_1_inst_00 : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => mulByte_1_inst_00_rhs,
    o   => mulByte_1_inst_00_o
  );
  mulByte_2_inst_02 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_02_rhs,
    o   => mulByte_2_inst_02_o
  );
  mulByte_2_inst_03 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_03_rhs,
    o   => mulByte_2_inst_03_o
  );
  mulByte_2_inst_04 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_04_rhs,
    o   => mulByte_2_inst_04_o
  );
  mulByte_0_inst_01 : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => mulByte_0_inst_01_rhs,
    o   => mulByte_0_inst_01_o
  );
  mulByte_1_inst_01 : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => mulByte_1_inst_01_rhs,
    o   => mulByte_1_inst_01_o
  );
  mulByte_1_inst_02 : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => mulByte_1_inst_02_rhs,
    o   => mulByte_1_inst_02_o
  );
  mulByte_2_inst_05 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_05_rhs,
    o   => mulByte_2_inst_05_o
  );
  mulByte_2_inst_06 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_06_rhs,
    o   => mulByte_2_inst_06_o
  );
  mulByte_0_inst_02 : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => mulByte_0_inst_02_rhs,
    o   => mulByte_0_inst_02_o
  );
  mulByte_0_inst_03 : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => mulByte_0_inst_03_rhs,
    o   => mulByte_0_inst_03_o
  );
  mulByte_1_inst_03 : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => mulByte_1_inst_03_rhs,
    o   => mulByte_1_inst_03_o
  );
  mulByte_2_inst_07 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_07_rhs,
    o   => mulByte_2_inst_07_o
  );
  mulByte_2_inst_08 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_08_rhs,
    o   => mulByte_2_inst_08_o
  );
  mulByte_2_inst_09 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_09_rhs,
    o   => mulByte_2_inst_09_o
  );
  mulByte_0_inst_04 : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => mulByte_0_inst_04_rhs,
    o   => mulByte_0_inst_04_o
  );
  mulByte_1_inst_04 : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => mulByte_1_inst_04_rhs,
    o   => mulByte_1_inst_04_o
  );
  mulByte_2_inst_10 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_10_rhs,
    o   => mulByte_2_inst_10_o
  );
  mulByte_2_inst_11 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_11_rhs,
    o   => mulByte_2_inst_11_o
  );
  mulByte_2_inst_12 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_12_rhs,
    o   => mulByte_2_inst_12_o
  );
  mulByte_0_inst_05 : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => mulByte_0_inst_05_rhs,
    o   => mulByte_0_inst_05_o
  );
  mulByte_1_inst_05 : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => mulByte_1_inst_05_rhs,
    o   => mulByte_1_inst_05_o
  );
  mulByte_1_inst_06 : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => mulByte_1_inst_06_rhs,
    o   => mulByte_1_inst_06_o
  );
  mulByte_2_inst_13 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_13_rhs,
    o   => mulByte_2_inst_13_o
  );
  mulByte_2_inst_14 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_14_rhs,
    o   => mulByte_2_inst_14_o
  );
  mulByte_0_inst_06 : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => mulByte_0_inst_06_rhs,
    o   => mulByte_0_inst_06_o
  );
  mulByte_0_inst_07 : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => mulByte_0_inst_07_rhs,
    o   => mulByte_0_inst_07_o
  );
  mulByte_1_inst_07 : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => mulByte_1_inst_07_rhs,
    o   => mulByte_1_inst_07_o
  );
  mulByte_2_inst_15 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_15_rhs,
    o   => mulByte_2_inst_15_o
  );
  mulByte_2_inst_16 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_16_rhs,
    o   => mulByte_2_inst_16_o
  );
  mulByte_2_inst_17 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_17_rhs,
    o   => mulByte_2_inst_17_o
  );
  mulByte_0_inst_08 : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => mulByte_0_inst_08_rhs,
    o   => mulByte_0_inst_08_o
  );
  mulByte_1_inst_08 : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => mulByte_1_inst_08_rhs,
    o   => mulByte_1_inst_08_o
  );
  mulByte_2_inst_18 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_18_rhs,
    o   => mulByte_2_inst_18_o
  );
  mulByte_2_inst_19 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_19_rhs,
    o   => mulByte_2_inst_19_o
  );
  mulByte_2_inst_20 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_20_rhs,
    o   => mulByte_2_inst_20_o
  );
  mulByte_0_inst_09 : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => mulByte_0_inst_09_rhs,
    o   => mulByte_0_inst_09_o
  );
  mulByte_1_inst_09 : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => mulByte_1_inst_09_rhs,
    o   => mulByte_1_inst_09_o
  );
  mulByte_1_inst_10 : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => mulByte_1_inst_10_rhs,
    o   => mulByte_1_inst_10_o
  );
  mulByte_2_inst_21 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_21_rhs,
    o   => mulByte_2_inst_21_o
  );
  mulByte_2_inst_22 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_22_rhs,
    o   => mulByte_2_inst_22_o
  );
  mulByte_0_inst_10 : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => mulByte_0_inst_10_rhs,
    o   => mulByte_0_inst_10_o
  );
  mulByte_0_inst_11 : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => mulByte_0_inst_11_rhs,
    o   => mulByte_0_inst_11_o
  );
  mulByte_1_inst_11 : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => mulByte_1_inst_11_rhs,
    o   => mulByte_1_inst_11_o
  );
  mulByte_2_inst_23 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_23_rhs,
    o   => mulByte_2_inst_23_o
  );
  mulByte_2_inst_24 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_24_rhs,
    o   => mulByte_2_inst_24_o
  );
  mulByte_2_inst_25 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_25_rhs,
    o   => mulByte_2_inst_25_o
  );
  mulByte_0_inst_12 : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => mulByte_0_inst_12_rhs,
    o   => mulByte_0_inst_12_o
  );
  mulByte_1_inst_12 : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => mulByte_1_inst_12_rhs,
    o   => mulByte_1_inst_12_o
  );
  mulByte_2_inst_26 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_26_rhs,
    o   => mulByte_2_inst_26_o
  );
  mulByte_2_inst_27 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_27_rhs,
    o   => mulByte_2_inst_27_o
  );
  mulByte_2_inst_28 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_28_rhs,
    o   => mulByte_2_inst_28_o
  );
  mulByte_0_inst_13 : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => mulByte_0_inst_13_rhs,
    o   => mulByte_0_inst_13_o
  );
  mulByte_1_inst_13 : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => mulByte_1_inst_13_rhs,
    o   => mulByte_1_inst_13_o
  );
  mulByte_1_inst_14 : entity work.mulByte_1(mulByte_1_arch) generic map (
    lhs => x"03"
  ) port map (
    rhs => mulByte_1_inst_14_rhs,
    o   => mulByte_1_inst_14_o
  );
  mulByte_2_inst_29 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_29_rhs,
    o   => mulByte_2_inst_29_o
  );
  mulByte_2_inst_30 : entity work.mulByte_2(mulByte_2_arch) generic map (
    lhs => x"01"
  ) port map (
    rhs => mulByte_2_inst_30_rhs,
    o   => mulByte_2_inst_30_o
  );
  mulByte_0_inst_14 : entity work.mulByte_0(mulByte_0_arch) generic map (
    lhs => x"02"
  ) port map (
    rhs => mulByte_0_inst_14_rhs,
    o   => mulByte_0_inst_14_o
  );
  o_part_mulByte_0_inst_rhs <= state(0)(0);
  o_part_mulByte_1_inst_rhs <= state(0)(1);
  o_part_mulByte_2_inst_rhs <= state(0)(2);
  mulByte_2_inst_00_rhs <= state(0)(3);
  mulByte_2_inst_01_rhs <= state(0)(0);
  mulByte_0_inst_00_rhs <= state(0)(1);
  mulByte_1_inst_00_rhs <= state(0)(2);
  mulByte_2_inst_02_rhs <= state(0)(3);
  mulByte_2_inst_03_rhs <= state(0)(0);
  mulByte_2_inst_04_rhs <= state(0)(1);
  mulByte_0_inst_01_rhs <= state(0)(2);
  mulByte_1_inst_01_rhs <= state(0)(3);
  mulByte_1_inst_02_rhs <= state(0)(0);
  mulByte_2_inst_05_rhs <= state(0)(1);
  mulByte_2_inst_06_rhs <= state(0)(2);
  mulByte_0_inst_02_rhs <= state(0)(3);
  mulByte_0_inst_03_rhs <= state(1)(0);
  mulByte_1_inst_03_rhs <= state(1)(1);
  mulByte_2_inst_07_rhs <= state(1)(2);
  mulByte_2_inst_08_rhs <= state(1)(3);
  mulByte_2_inst_09_rhs <= state(1)(0);
  mulByte_0_inst_04_rhs <= state(1)(1);
  mulByte_1_inst_04_rhs <= state(1)(2);
  mulByte_2_inst_10_rhs <= state(1)(3);
  mulByte_2_inst_11_rhs <= state(1)(0);
  mulByte_2_inst_12_rhs <= state(1)(1);
  mulByte_0_inst_05_rhs <= state(1)(2);
  mulByte_1_inst_05_rhs <= state(1)(3);
  mulByte_1_inst_06_rhs <= state(1)(0);
  mulByte_2_inst_13_rhs <= state(1)(1);
  mulByte_2_inst_14_rhs <= state(1)(2);
  mulByte_0_inst_06_rhs <= state(1)(3);
  mulByte_0_inst_07_rhs <= state(2)(0);
  mulByte_1_inst_07_rhs <= state(2)(1);
  mulByte_2_inst_15_rhs <= state(2)(2);
  mulByte_2_inst_16_rhs <= state(2)(3);
  mulByte_2_inst_17_rhs <= state(2)(0);
  mulByte_0_inst_08_rhs <= state(2)(1);
  mulByte_1_inst_08_rhs <= state(2)(2);
  mulByte_2_inst_18_rhs <= state(2)(3);
  mulByte_2_inst_19_rhs <= state(2)(0);
  mulByte_2_inst_20_rhs <= state(2)(1);
  mulByte_0_inst_09_rhs <= state(2)(2);
  mulByte_1_inst_09_rhs <= state(2)(3);
  mulByte_1_inst_10_rhs <= state(2)(0);
  mulByte_2_inst_21_rhs <= state(2)(1);
  mulByte_2_inst_22_rhs <= state(2)(2);
  mulByte_0_inst_10_rhs <= state(2)(3);
  mulByte_0_inst_11_rhs <= state(3)(0);
  mulByte_1_inst_11_rhs <= state(3)(1);
  mulByte_2_inst_23_rhs <= state(3)(2);
  mulByte_2_inst_24_rhs <= state(3)(3);
  mulByte_2_inst_25_rhs <= state(3)(0);
  mulByte_0_inst_12_rhs <= state(3)(1);
  mulByte_1_inst_12_rhs <= state(3)(2);
  mulByte_2_inst_26_rhs <= state(3)(3);
  mulByte_2_inst_27_rhs <= state(3)(0);
  mulByte_2_inst_28_rhs <= state(3)(1);
  mulByte_0_inst_13_rhs <= state(3)(2);
  mulByte_1_inst_13_rhs <= state(3)(3);
  mulByte_1_inst_14_rhs <= state(3)(0);
  mulByte_2_inst_29_rhs <= state(3)(1);
  mulByte_2_inst_30_rhs <= state(3)(2);
  mulByte_0_inst_14_rhs <= state(3)(3);
  o     <= (
    0   => (
      0 => ((o_part_mulByte_0_inst_o xor o_part_mulByte_1_inst_o) xor o_part_mulByte_2_inst_o) xor mulByte_2_inst_00_o,
      1 => ((mulByte_2_inst_01_o xor mulByte_0_inst_00_o) xor mulByte_1_inst_00_o) xor mulByte_2_inst_02_o,
      2 => ((mulByte_2_inst_03_o xor mulByte_2_inst_04_o) xor mulByte_0_inst_01_o) xor mulByte_1_inst_01_o,
      3 => ((mulByte_1_inst_02_o xor mulByte_2_inst_05_o) xor mulByte_2_inst_06_o) xor mulByte_0_inst_02_o
    ),
    1   => (
      0 => ((mulByte_0_inst_03_o xor mulByte_1_inst_03_o) xor mulByte_2_inst_07_o) xor mulByte_2_inst_08_o,
      1 => ((mulByte_2_inst_09_o xor mulByte_0_inst_04_o) xor mulByte_1_inst_04_o) xor mulByte_2_inst_10_o,
      2 => ((mulByte_2_inst_11_o xor mulByte_2_inst_12_o) xor mulByte_0_inst_05_o) xor mulByte_1_inst_05_o,
      3 => ((mulByte_1_inst_06_o xor mulByte_2_inst_13_o) xor mulByte_2_inst_14_o) xor mulByte_0_inst_06_o
    ),
    2   => (
      0 => ((mulByte_0_inst_07_o xor mulByte_1_inst_07_o) xor mulByte_2_inst_15_o) xor mulByte_2_inst_16_o,
      1 => ((mulByte_2_inst_17_o xor mulByte_0_inst_08_o) xor mulByte_1_inst_08_o) xor mulByte_2_inst_18_o,
      2 => ((mulByte_2_inst_19_o xor mulByte_2_inst_20_o) xor mulByte_0_inst_09_o) xor mulByte_1_inst_09_o,
      3 => ((mulByte_1_inst_10_o xor mulByte_2_inst_21_o) xor mulByte_2_inst_22_o) xor mulByte_0_inst_10_o
    ),
    3   => (
      0 => ((mulByte_0_inst_11_o xor mulByte_1_inst_11_o) xor mulByte_2_inst_23_o) xor mulByte_2_inst_24_o,
      1 => ((mulByte_2_inst_25_o xor mulByte_0_inst_12_o) xor mulByte_1_inst_12_o) xor mulByte_2_inst_26_o,
      2 => ((mulByte_2_inst_27_o xor mulByte_2_inst_28_o) xor mulByte_0_inst_13_o) xor mulByte_1_inst_13_o,
      3 => ((mulByte_1_inst_14_o xor mulByte_2_inst_29_o) xor mulByte_2_inst_30_o) xor mulByte_0_inst_14_o
    )
  );
end mixColumns_arch;
