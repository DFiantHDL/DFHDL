`ifndef BLINKER_DEFS
`define BLINKER_DEFS
`endif
`ifndef BLINKER_DEFS_MODULE
`define BLINKER_DEFS_MODULE
`else

`undef BLINKER_DEFS_MODULE
`endif

