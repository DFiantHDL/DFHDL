`ifndef TRUEDPR_DEFS
`define TRUEDPR_DEFS

`endif
