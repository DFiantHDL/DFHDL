library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.dfhdl_pkg.all;

package LeftShift2_pkg is
end package LeftShift2_pkg;

package body LeftShift2_pkg is
end package body LeftShift2_pkg;
