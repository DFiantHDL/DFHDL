library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.dfhdl_pkg.all;

package RegFile_pkg is
end package RegFile_pkg;

package body RegFile_pkg is
end package body RegFile_pkg;
