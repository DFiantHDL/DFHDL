`ifndef COUNTER_DEFS
`define COUNTER_DEFS

`endif
`ifndef COUNTER_DEFS_MODULE
`define COUNTER_DEFS_MODULE
`else

`undef COUNTER_DEFS_MODULE
`endif

