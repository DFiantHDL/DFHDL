`ifndef LEFTSHIFT2_DEFS
`define LEFTSHIFT2_DEFS

`endif
`ifndef LEFTSHIFT2_DEFS_MODULE
`define LEFTSHIFT2_DEFS_MODULE
`else

`undef LEFTSHIFT2_DEFS_MODULE
`endif

