`ifndef FULLADDERN_DEFS
`define FULLADDERN_DEFS

`endif
`ifndef FULLADDERN_DEFS_MODULE
`define FULLADDERN_DEFS_MODULE
`else

`undef FULLADDERN_DEFS_MODULE
`endif

