library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.dfhdl_pkg.all;

package FullAdderN_pkg is

end package FullAdderN_pkg;

package body FullAdderN_pkg is

end package body FullAdderN_pkg;
