`default_nettype none
`timescale 1ns/1ps
`include "CipherNoOpaques_defs.vh"

module sbox(
  lhs,
  o
);
  `include "dfhdl_defs.vh"
  `include "CipherNoOpaques_defs.vh"
  `sboxLookupTable_def
  input  wire  [7:0] lhs;
  output wire [7:0]  o;
  reg [7:0] sboxLookupTable_rom [0:255];
  initial begin : sboxLookupTable_rom_init
    sboxLookupTable_rom[0]   = sboxLookupTable[2047:2040];
    sboxLookupTable_rom[1]   = sboxLookupTable[2039:2032];
    sboxLookupTable_rom[2]   = sboxLookupTable[2031:2024];
    sboxLookupTable_rom[3]   = sboxLookupTable[2023:2016];
    sboxLookupTable_rom[4]   = sboxLookupTable[2015:2008];
    sboxLookupTable_rom[5]   = sboxLookupTable[2007:2000];
    sboxLookupTable_rom[6]   = sboxLookupTable[1999:1992];
    sboxLookupTable_rom[7]   = sboxLookupTable[1991:1984];
    sboxLookupTable_rom[8]   = sboxLookupTable[1983:1976];
    sboxLookupTable_rom[9]   = sboxLookupTable[1975:1968];
    sboxLookupTable_rom[10]  = sboxLookupTable[1967:1960];
    sboxLookupTable_rom[11]  = sboxLookupTable[1959:1952];
    sboxLookupTable_rom[12]  = sboxLookupTable[1951:1944];
    sboxLookupTable_rom[13]  = sboxLookupTable[1943:1936];
    sboxLookupTable_rom[14]  = sboxLookupTable[1935:1928];
    sboxLookupTable_rom[15]  = sboxLookupTable[1927:1920];
    sboxLookupTable_rom[16]  = sboxLookupTable[1919:1912];
    sboxLookupTable_rom[17]  = sboxLookupTable[1911:1904];
    sboxLookupTable_rom[18]  = sboxLookupTable[1903:1896];
    sboxLookupTable_rom[19]  = sboxLookupTable[1895:1888];
    sboxLookupTable_rom[20]  = sboxLookupTable[1887:1880];
    sboxLookupTable_rom[21]  = sboxLookupTable[1879:1872];
    sboxLookupTable_rom[22]  = sboxLookupTable[1871:1864];
    sboxLookupTable_rom[23]  = sboxLookupTable[1863:1856];
    sboxLookupTable_rom[24]  = sboxLookupTable[1855:1848];
    sboxLookupTable_rom[25]  = sboxLookupTable[1847:1840];
    sboxLookupTable_rom[26]  = sboxLookupTable[1839:1832];
    sboxLookupTable_rom[27]  = sboxLookupTable[1831:1824];
    sboxLookupTable_rom[28]  = sboxLookupTable[1823:1816];
    sboxLookupTable_rom[29]  = sboxLookupTable[1815:1808];
    sboxLookupTable_rom[30]  = sboxLookupTable[1807:1800];
    sboxLookupTable_rom[31]  = sboxLookupTable[1799:1792];
    sboxLookupTable_rom[32]  = sboxLookupTable[1791:1784];
    sboxLookupTable_rom[33]  = sboxLookupTable[1783:1776];
    sboxLookupTable_rom[34]  = sboxLookupTable[1775:1768];
    sboxLookupTable_rom[35]  = sboxLookupTable[1767:1760];
    sboxLookupTable_rom[36]  = sboxLookupTable[1759:1752];
    sboxLookupTable_rom[37]  = sboxLookupTable[1751:1744];
    sboxLookupTable_rom[38]  = sboxLookupTable[1743:1736];
    sboxLookupTable_rom[39]  = sboxLookupTable[1735:1728];
    sboxLookupTable_rom[40]  = sboxLookupTable[1727:1720];
    sboxLookupTable_rom[41]  = sboxLookupTable[1719:1712];
    sboxLookupTable_rom[42]  = sboxLookupTable[1711:1704];
    sboxLookupTable_rom[43]  = sboxLookupTable[1703:1696];
    sboxLookupTable_rom[44]  = sboxLookupTable[1695:1688];
    sboxLookupTable_rom[45]  = sboxLookupTable[1687:1680];
    sboxLookupTable_rom[46]  = sboxLookupTable[1679:1672];
    sboxLookupTable_rom[47]  = sboxLookupTable[1671:1664];
    sboxLookupTable_rom[48]  = sboxLookupTable[1663:1656];
    sboxLookupTable_rom[49]  = sboxLookupTable[1655:1648];
    sboxLookupTable_rom[50]  = sboxLookupTable[1647:1640];
    sboxLookupTable_rom[51]  = sboxLookupTable[1639:1632];
    sboxLookupTable_rom[52]  = sboxLookupTable[1631:1624];
    sboxLookupTable_rom[53]  = sboxLookupTable[1623:1616];
    sboxLookupTable_rom[54]  = sboxLookupTable[1615:1608];
    sboxLookupTable_rom[55]  = sboxLookupTable[1607:1600];
    sboxLookupTable_rom[56]  = sboxLookupTable[1599:1592];
    sboxLookupTable_rom[57]  = sboxLookupTable[1591:1584];
    sboxLookupTable_rom[58]  = sboxLookupTable[1583:1576];
    sboxLookupTable_rom[59]  = sboxLookupTable[1575:1568];
    sboxLookupTable_rom[60]  = sboxLookupTable[1567:1560];
    sboxLookupTable_rom[61]  = sboxLookupTable[1559:1552];
    sboxLookupTable_rom[62]  = sboxLookupTable[1551:1544];
    sboxLookupTable_rom[63]  = sboxLookupTable[1543:1536];
    sboxLookupTable_rom[64]  = sboxLookupTable[1535:1528];
    sboxLookupTable_rom[65]  = sboxLookupTable[1527:1520];
    sboxLookupTable_rom[66]  = sboxLookupTable[1519:1512];
    sboxLookupTable_rom[67]  = sboxLookupTable[1511:1504];
    sboxLookupTable_rom[68]  = sboxLookupTable[1503:1496];
    sboxLookupTable_rom[69]  = sboxLookupTable[1495:1488];
    sboxLookupTable_rom[70]  = sboxLookupTable[1487:1480];
    sboxLookupTable_rom[71]  = sboxLookupTable[1479:1472];
    sboxLookupTable_rom[72]  = sboxLookupTable[1471:1464];
    sboxLookupTable_rom[73]  = sboxLookupTable[1463:1456];
    sboxLookupTable_rom[74]  = sboxLookupTable[1455:1448];
    sboxLookupTable_rom[75]  = sboxLookupTable[1447:1440];
    sboxLookupTable_rom[76]  = sboxLookupTable[1439:1432];
    sboxLookupTable_rom[77]  = sboxLookupTable[1431:1424];
    sboxLookupTable_rom[78]  = sboxLookupTable[1423:1416];
    sboxLookupTable_rom[79]  = sboxLookupTable[1415:1408];
    sboxLookupTable_rom[80]  = sboxLookupTable[1407:1400];
    sboxLookupTable_rom[81]  = sboxLookupTable[1399:1392];
    sboxLookupTable_rom[82]  = sboxLookupTable[1391:1384];
    sboxLookupTable_rom[83]  = sboxLookupTable[1383:1376];
    sboxLookupTable_rom[84]  = sboxLookupTable[1375:1368];
    sboxLookupTable_rom[85]  = sboxLookupTable[1367:1360];
    sboxLookupTable_rom[86]  = sboxLookupTable[1359:1352];
    sboxLookupTable_rom[87]  = sboxLookupTable[1351:1344];
    sboxLookupTable_rom[88]  = sboxLookupTable[1343:1336];
    sboxLookupTable_rom[89]  = sboxLookupTable[1335:1328];
    sboxLookupTable_rom[90]  = sboxLookupTable[1327:1320];
    sboxLookupTable_rom[91]  = sboxLookupTable[1319:1312];
    sboxLookupTable_rom[92]  = sboxLookupTable[1311:1304];
    sboxLookupTable_rom[93]  = sboxLookupTable[1303:1296];
    sboxLookupTable_rom[94]  = sboxLookupTable[1295:1288];
    sboxLookupTable_rom[95]  = sboxLookupTable[1287:1280];
    sboxLookupTable_rom[96]  = sboxLookupTable[1279:1272];
    sboxLookupTable_rom[97]  = sboxLookupTable[1271:1264];
    sboxLookupTable_rom[98]  = sboxLookupTable[1263:1256];
    sboxLookupTable_rom[99]  = sboxLookupTable[1255:1248];
    sboxLookupTable_rom[100] = sboxLookupTable[1247:1240];
    sboxLookupTable_rom[101] = sboxLookupTable[1239:1232];
    sboxLookupTable_rom[102] = sboxLookupTable[1231:1224];
    sboxLookupTable_rom[103] = sboxLookupTable[1223:1216];
    sboxLookupTable_rom[104] = sboxLookupTable[1215:1208];
    sboxLookupTable_rom[105] = sboxLookupTable[1207:1200];
    sboxLookupTable_rom[106] = sboxLookupTable[1199:1192];
    sboxLookupTable_rom[107] = sboxLookupTable[1191:1184];
    sboxLookupTable_rom[108] = sboxLookupTable[1183:1176];
    sboxLookupTable_rom[109] = sboxLookupTable[1175:1168];
    sboxLookupTable_rom[110] = sboxLookupTable[1167:1160];
    sboxLookupTable_rom[111] = sboxLookupTable[1159:1152];
    sboxLookupTable_rom[112] = sboxLookupTable[1151:1144];
    sboxLookupTable_rom[113] = sboxLookupTable[1143:1136];
    sboxLookupTable_rom[114] = sboxLookupTable[1135:1128];
    sboxLookupTable_rom[115] = sboxLookupTable[1127:1120];
    sboxLookupTable_rom[116] = sboxLookupTable[1119:1112];
    sboxLookupTable_rom[117] = sboxLookupTable[1111:1104];
    sboxLookupTable_rom[118] = sboxLookupTable[1103:1096];
    sboxLookupTable_rom[119] = sboxLookupTable[1095:1088];
    sboxLookupTable_rom[120] = sboxLookupTable[1087:1080];
    sboxLookupTable_rom[121] = sboxLookupTable[1079:1072];
    sboxLookupTable_rom[122] = sboxLookupTable[1071:1064];
    sboxLookupTable_rom[123] = sboxLookupTable[1063:1056];
    sboxLookupTable_rom[124] = sboxLookupTable[1055:1048];
    sboxLookupTable_rom[125] = sboxLookupTable[1047:1040];
    sboxLookupTable_rom[126] = sboxLookupTable[1039:1032];
    sboxLookupTable_rom[127] = sboxLookupTable[1031:1024];
    sboxLookupTable_rom[128] = sboxLookupTable[1023:1016];
    sboxLookupTable_rom[129] = sboxLookupTable[1015:1008];
    sboxLookupTable_rom[130] = sboxLookupTable[1007:1000];
    sboxLookupTable_rom[131] = sboxLookupTable[999:992];
    sboxLookupTable_rom[132] = sboxLookupTable[991:984];
    sboxLookupTable_rom[133] = sboxLookupTable[983:976];
    sboxLookupTable_rom[134] = sboxLookupTable[975:968];
    sboxLookupTable_rom[135] = sboxLookupTable[967:960];
    sboxLookupTable_rom[136] = sboxLookupTable[959:952];
    sboxLookupTable_rom[137] = sboxLookupTable[951:944];
    sboxLookupTable_rom[138] = sboxLookupTable[943:936];
    sboxLookupTable_rom[139] = sboxLookupTable[935:928];
    sboxLookupTable_rom[140] = sboxLookupTable[927:920];
    sboxLookupTable_rom[141] = sboxLookupTable[919:912];
    sboxLookupTable_rom[142] = sboxLookupTable[911:904];
    sboxLookupTable_rom[143] = sboxLookupTable[903:896];
    sboxLookupTable_rom[144] = sboxLookupTable[895:888];
    sboxLookupTable_rom[145] = sboxLookupTable[887:880];
    sboxLookupTable_rom[146] = sboxLookupTable[879:872];
    sboxLookupTable_rom[147] = sboxLookupTable[871:864];
    sboxLookupTable_rom[148] = sboxLookupTable[863:856];
    sboxLookupTable_rom[149] = sboxLookupTable[855:848];
    sboxLookupTable_rom[150] = sboxLookupTable[847:840];
    sboxLookupTable_rom[151] = sboxLookupTable[839:832];
    sboxLookupTable_rom[152] = sboxLookupTable[831:824];
    sboxLookupTable_rom[153] = sboxLookupTable[823:816];
    sboxLookupTable_rom[154] = sboxLookupTable[815:808];
    sboxLookupTable_rom[155] = sboxLookupTable[807:800];
    sboxLookupTable_rom[156] = sboxLookupTable[799:792];
    sboxLookupTable_rom[157] = sboxLookupTable[791:784];
    sboxLookupTable_rom[158] = sboxLookupTable[783:776];
    sboxLookupTable_rom[159] = sboxLookupTable[775:768];
    sboxLookupTable_rom[160] = sboxLookupTable[767:760];
    sboxLookupTable_rom[161] = sboxLookupTable[759:752];
    sboxLookupTable_rom[162] = sboxLookupTable[751:744];
    sboxLookupTable_rom[163] = sboxLookupTable[743:736];
    sboxLookupTable_rom[164] = sboxLookupTable[735:728];
    sboxLookupTable_rom[165] = sboxLookupTable[727:720];
    sboxLookupTable_rom[166] = sboxLookupTable[719:712];
    sboxLookupTable_rom[167] = sboxLookupTable[711:704];
    sboxLookupTable_rom[168] = sboxLookupTable[703:696];
    sboxLookupTable_rom[169] = sboxLookupTable[695:688];
    sboxLookupTable_rom[170] = sboxLookupTable[687:680];
    sboxLookupTable_rom[171] = sboxLookupTable[679:672];
    sboxLookupTable_rom[172] = sboxLookupTable[671:664];
    sboxLookupTable_rom[173] = sboxLookupTable[663:656];
    sboxLookupTable_rom[174] = sboxLookupTable[655:648];
    sboxLookupTable_rom[175] = sboxLookupTable[647:640];
    sboxLookupTable_rom[176] = sboxLookupTable[639:632];
    sboxLookupTable_rom[177] = sboxLookupTable[631:624];
    sboxLookupTable_rom[178] = sboxLookupTable[623:616];
    sboxLookupTable_rom[179] = sboxLookupTable[615:608];
    sboxLookupTable_rom[180] = sboxLookupTable[607:600];
    sboxLookupTable_rom[181] = sboxLookupTable[599:592];
    sboxLookupTable_rom[182] = sboxLookupTable[591:584];
    sboxLookupTable_rom[183] = sboxLookupTable[583:576];
    sboxLookupTable_rom[184] = sboxLookupTable[575:568];
    sboxLookupTable_rom[185] = sboxLookupTable[567:560];
    sboxLookupTable_rom[186] = sboxLookupTable[559:552];
    sboxLookupTable_rom[187] = sboxLookupTable[551:544];
    sboxLookupTable_rom[188] = sboxLookupTable[543:536];
    sboxLookupTable_rom[189] = sboxLookupTable[535:528];
    sboxLookupTable_rom[190] = sboxLookupTable[527:520];
    sboxLookupTable_rom[191] = sboxLookupTable[519:512];
    sboxLookupTable_rom[192] = sboxLookupTable[511:504];
    sboxLookupTable_rom[193] = sboxLookupTable[503:496];
    sboxLookupTable_rom[194] = sboxLookupTable[495:488];
    sboxLookupTable_rom[195] = sboxLookupTable[487:480];
    sboxLookupTable_rom[196] = sboxLookupTable[479:472];
    sboxLookupTable_rom[197] = sboxLookupTable[471:464];
    sboxLookupTable_rom[198] = sboxLookupTable[463:456];
    sboxLookupTable_rom[199] = sboxLookupTable[455:448];
    sboxLookupTable_rom[200] = sboxLookupTable[447:440];
    sboxLookupTable_rom[201] = sboxLookupTable[439:432];
    sboxLookupTable_rom[202] = sboxLookupTable[431:424];
    sboxLookupTable_rom[203] = sboxLookupTable[423:416];
    sboxLookupTable_rom[204] = sboxLookupTable[415:408];
    sboxLookupTable_rom[205] = sboxLookupTable[407:400];
    sboxLookupTable_rom[206] = sboxLookupTable[399:392];
    sboxLookupTable_rom[207] = sboxLookupTable[391:384];
    sboxLookupTable_rom[208] = sboxLookupTable[383:376];
    sboxLookupTable_rom[209] = sboxLookupTable[375:368];
    sboxLookupTable_rom[210] = sboxLookupTable[367:360];
    sboxLookupTable_rom[211] = sboxLookupTable[359:352];
    sboxLookupTable_rom[212] = sboxLookupTable[351:344];
    sboxLookupTable_rom[213] = sboxLookupTable[343:336];
    sboxLookupTable_rom[214] = sboxLookupTable[335:328];
    sboxLookupTable_rom[215] = sboxLookupTable[327:320];
    sboxLookupTable_rom[216] = sboxLookupTable[319:312];
    sboxLookupTable_rom[217] = sboxLookupTable[311:304];
    sboxLookupTable_rom[218] = sboxLookupTable[303:296];
    sboxLookupTable_rom[219] = sboxLookupTable[295:288];
    sboxLookupTable_rom[220] = sboxLookupTable[287:280];
    sboxLookupTable_rom[221] = sboxLookupTable[279:272];
    sboxLookupTable_rom[222] = sboxLookupTable[271:264];
    sboxLookupTable_rom[223] = sboxLookupTable[263:256];
    sboxLookupTable_rom[224] = sboxLookupTable[255:248];
    sboxLookupTable_rom[225] = sboxLookupTable[247:240];
    sboxLookupTable_rom[226] = sboxLookupTable[239:232];
    sboxLookupTable_rom[227] = sboxLookupTable[231:224];
    sboxLookupTable_rom[228] = sboxLookupTable[223:216];
    sboxLookupTable_rom[229] = sboxLookupTable[215:208];
    sboxLookupTable_rom[230] = sboxLookupTable[207:200];
    sboxLookupTable_rom[231] = sboxLookupTable[199:192];
    sboxLookupTable_rom[232] = sboxLookupTable[191:184];
    sboxLookupTable_rom[233] = sboxLookupTable[183:176];
    sboxLookupTable_rom[234] = sboxLookupTable[175:168];
    sboxLookupTable_rom[235] = sboxLookupTable[167:160];
    sboxLookupTable_rom[236] = sboxLookupTable[159:152];
    sboxLookupTable_rom[237] = sboxLookupTable[151:144];
    sboxLookupTable_rom[238] = sboxLookupTable[143:136];
    sboxLookupTable_rom[239] = sboxLookupTable[135:128];
    sboxLookupTable_rom[240] = sboxLookupTable[127:120];
    sboxLookupTable_rom[241] = sboxLookupTable[119:112];
    sboxLookupTable_rom[242] = sboxLookupTable[111:104];
    sboxLookupTable_rom[243] = sboxLookupTable[103:96];
    sboxLookupTable_rom[244] = sboxLookupTable[95:88];
    sboxLookupTable_rom[245] = sboxLookupTable[87:80];
    sboxLookupTable_rom[246] = sboxLookupTable[79:72];
    sboxLookupTable_rom[247] = sboxLookupTable[71:64];
    sboxLookupTable_rom[248] = sboxLookupTable[63:56];
    sboxLookupTable_rom[249] = sboxLookupTable[55:48];
    sboxLookupTable_rom[250] = sboxLookupTable[47:40];
    sboxLookupTable_rom[251] = sboxLookupTable[39:32];
    sboxLookupTable_rom[252] = sboxLookupTable[31:24];
    sboxLookupTable_rom[253] = sboxLookupTable[23:16];
    sboxLookupTable_rom[254] = sboxLookupTable[15:8];
    sboxLookupTable_rom[255] = sboxLookupTable[7:0];
  end
  assign o = sboxLookupTable_rom[lhs];
endmodule
