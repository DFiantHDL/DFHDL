`ifndef TRUEDPR_DEFS
`define TRUEDPR_DEFS
`endif
`ifndef TRUEDPR_DEFS_MODULE
`define TRUEDPR_DEFS_MODULE
`else

`undef TRUEDPR_DEFS_MODULE
`endif

