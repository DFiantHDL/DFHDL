`ifndef COUNTER_DEFS
`define COUNTER_DEFS
`endif
