`ifndef BLINKER_DEFS
`define BLINKER_DEFS
`endif
