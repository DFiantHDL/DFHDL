library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.dfhdl_pkg.all;

package LeftShiftBasic_pkg is

end package LeftShiftBasic_pkg;

package body LeftShiftBasic_pkg is

end package body LeftShiftBasic_pkg;
