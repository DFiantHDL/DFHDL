library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.dfhdl_pkg.all;

package LeftShiftGen_pkg is

end package LeftShiftGen_pkg;

package body LeftShiftGen_pkg is

end package body LeftShiftGen_pkg;
