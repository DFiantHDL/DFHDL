library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.dfhdl_pkg.all;

package Blinker_pkg is
end package Blinker_pkg;

package body Blinker_pkg is
end package body Blinker_pkg;
